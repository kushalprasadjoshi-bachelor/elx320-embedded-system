----------------------------------------------------------------------------------
-- Module Name:    Exp02_FullAdder - Behavioral 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Exp02_FullAdder is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           Cin : in  STD_LOGIC;
           Sum : out  STD_LOGIC;
           Cout : out  STD_LOGIC);
end Exp02_FullAdder;

architecture Behavioral of Exp02_FullAdder is

begin
    -- Sum is the XOR of A, B, and Cin
    Sum <= A XOR B XOR Cin;
    
    -- Carry output is generated by:
    -- (A AND B) OR (B AND Cin) OR (A AND Cin)
    Cout <= (A AND B) OR (B AND Cin) OR (A AND Cin);

end Behavioral;

