----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:30:58 01/21/2026 
-- Design Name: 
-- Module Name:    Exp02_FullAdder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Exp02_FullAdder is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           Cin : in  STD_LOGIC;
           Sum : out  STD_LOGIC;
           Cout : out  STD_LOGIC);
end Exp02_FullAdder;

architecture Behavioral of Exp02_FullAdder is

begin
    -- Sum is the XOR of A, B, and Cin
    Sum <= A XOR B XOR Cin;
    
    -- Carry output is generated by:
    -- (A AND B) OR (B AND Cin) OR (A AND Cin)
    Cout <= (A AND B) OR (B AND Cin) OR (A AND Cin);

end Behavioral;

